`include "adder.v"
`include "data_memory.v"
`include "memory_instruction.v"
`include "pc_ver.v"
`include "ALU.v"
`include "Register_files.v"
`include "risc_v_basic.v"


